------------------------------------------------------------------------------
--! Copyright (C) 2009 , Olivier Girard
--
--! Redistribution and use in source and binary forms, with or without
--! modification, are permitted provided that the following conditions
--! are met:
--!     * Redistributions of source code must retain the above copyright
--!       notice, this list of conditions and the following disclaimer.
--!     * Redistributions in binary form must reproduce the above copyright
--!       notice, this list of conditions and the following disclaimer in the
--!       documentation and/or other materials provided with the distribution.
--!     * Neither the name of the authors nor the names of its contributors
--!       may be used to endorse or promote products derived from this software
--!       without specific prior written permission.
--
--! THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
--! AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
--! IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
--! ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
--! LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--! OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
--! SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
--! INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
--! CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
--! ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF
--! THE POSSIBILITY OF SUCH DAMAGE
--
------------------------------------------------------------------------------
--
--! @file fmsp_clock_gate.vhd
--! 
--! @brief fpgaMSP430 Generic clock gate cell
--
--! @author Olivier Girard,    olgirard@gmail.com
--! @author Emmanuel Amadio,   emmanuel.amadio@gmail.com (VHDL Rewrite)
--
------------------------------------------------------------------------------
--! @version 1
--! @date: 2017-04-21
------------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;	--! standard unresolved logic UX01ZWLH-

entity fmsp_clock_gate is 
port (
	--! INPUTs
	clk			: in	std_logic;	--! Clock
	enable		: in	std_logic;	--! Clock enable
	scan_enable	: in	std_logic;	--! Scan enable (active during scan shifting)
	--! OUTPUTs
	gclk			: out	std_logic	--! Gated clock
);
end entity fmsp_clock_gate;

architecture RTL of fmsp_clock_gate is 

	signal	enable_in		: std_logic;
	signal	enable_latch	: std_logic;

begin
	
--=============================================================================
--! CLOCK GATE: LATCH + AND
--=============================================================================

--! Enable clock gate during scan shift
--! (the gate itself is checked with the scan capture cycle)
	enable_in	<= enable or scan_enable;

--! LATCH the enable signal
	LATCH_REG : process(clk,enable_in)
	begin
		if (not(clk) = '1') then
			enable_latch <= enable_in;
		end if;
	end process LATCH_REG;

	--! AND gate
	gclk <= clk and enable_latch;

end RTL; --! fmsp_clock_gate


